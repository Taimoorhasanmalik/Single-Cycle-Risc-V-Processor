module instr_mem_tb ();
    logic [31:0] addr,pc;
    instr_mem mem(pc,addr);
    initial begin
        pc = 0;
        #10;
        pc = 4;
        #10;
        pc = 8;
        #10;
        pc = 12;
        #10;
        pc = 16;
        #10;
        pc = 20;
        #10;
        pc = 24;
        #10;
        pc = 28;
        #10;
        pc = 32;
        #10;
        pc = 36;
        #10;
        pc = 40;
        #10;
        pc = 44;
        #10;
        pc = 48;
        #10;
        pc = 52;
        #10;
        pc = 56;
        #10;
        pc = 60;
        #10;
        pc = 64;
        #10;
        pc = 68;
        #10;
        pc = 72;
        #10;
        pc = 76;
        #10;
        pc = 80;
        #10;
        pc = 84;
        #10;
        pc = 88;
        #10;
        pc = 92;
        #10;
        pc = 96;
        #10;
        pc = 10;
        #10;
        pc = 104;
        #10;
        pc = 108;
        #10;
        pc = 112;
        #10;
        pc = 116;
        #10;
        pc = 120;
        #10;
        pc = 124;
        #10;
        pc = 128;
        #10;
        pc = 132;
        #10;
        pc = 136;
        #10;
        pc = 140;
        #10;
        pc = 144;
        #10;
        pc = 148;
        #10;
        pc = 152;
        #10;
        pc = 156;
        #10;
        pc = 160;
        #10;
        pc = 164;
        #10;
        pc = 168;
        #10;
        pc = 172;
        #10;
        pc = 176;
        #10;
        pc = 180;
        #10;
        pc = 184;
        #10;
        pc = 188;
        #10;
        pc = 192;
        #10;
        pc = 196;

    end


endmodule